module vga(
	input CLOCK_50,
	input rst,
	output hsync,
	output vsync	
);
	
endmodule